module	asyn_fifo#(
    parameter WIDTH = 8,
    parameter DEPTH = 16
)(
    input wclk,
    input rclk,
    input wrstn,
    input rrstn,
    input winc,
    input rinc,
    input [WIDTH-1:0] wdata,

    output wire wfull,
    output wire rempty,
    output wire [WIDTH-1:0] rdata
);

    // Internal signal definitions
    reg [$clog2(DEPTH):0] waddr, raddr;
    wire [$clog2(DEPTH):0] waddr_bin, raddr_bin;
    reg [$clog2(DEPTH):0] waddr_gray, raddr_gray;
    reg [$clog2(DEPTH):0] wptr, rptr;
    reg [$clog2(DEPTH):0] wptr_buff1, wptr_buff2, rptr_buff1, rptr_buff2;
    wire [$clog2(DEPTH):0] wptr_bin, rptr_bin;

    // Module instantiation
    dual_port_RAM #(.DEPTH(DEPTH), .WIDTH(WIDTH)) RAM(
        .wclk(wclk),
        .wenc(winc),
        .waddr(waddr_bin),
        .wdata(wdata),
        .rclk(rclk),
        .renc(rinc),
        .raddr(raddr_bin),
        .rdata(rdata)
    );

    // Pointer increment
    always @(posedge wclk or negedge wrstn) begin
        if (~wrstn)
            waddr <= 0;
        else if (winc && !wfull)
            waddr <= waddr + 1;
    end

    always @(posedge rclk or negedge rrstn) begin
        if (~rrstn)
            raddr <= 0;
        else if (rinc && !rempty)
            raddr <= raddr + 1;
    end

    // Convert to Gray code
    always @(waddr)
        waddr_gray <= waddr ^ (waddr >> 1);

    always @(raddr)
        raddr_gray <= raddr ^ (raddr >> 1);

    // Synchronize pointers
    always @(posedge wclk or negedge wrstn) begin
        if (~wrstn)
            wptr <= 0;
        else
            wptr <= waddr_gray;
    end

    always @(posedge rclk or negedge rrstn) begin
        if (~rrstn)
            rptr <= 0;
        else
            rptr <= raddr_gray;
    end

    // FIFO full and empty flags
    assign wfull = (wptr == (~rptr[WIDTH] & {rptr[WIDTH-1:0], 1'b1}));
    assign rempty = (wptr == rptr);

    // Binary address for RAM
    assign waddr_bin = waddr[WIDTH-1:0];
    assign raddr_bin = raddr[WIDTH-1:0];

endmodule
