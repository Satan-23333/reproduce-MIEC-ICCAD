module	dual_port_RAM #(
    parameter DEPTH = 16,
    parameter WIDTH = 8
)(
    input wclk,
    input rclk,
    input wenc,
    input [$clog2(DEPTH)-1:0] waddr,
    input [WIDTH-1:0] wdata,
    input renc,
    input [$clog2(DEPTH)-1:0] raddr,
    output reg [WIDTH-1:0] rdata
);
    reg [WIDTH-1:0] RAM_MEM [0:DEPTH-1];
    
    always @(posedge wclk)
        if(wenc)
            RAM_MEM[waddr] <= wdata;

    always @(posedge rclk)
        if(renc)
            rdata <= RAM_MEM[raddr];
endmodule
module	asyn_fifo#(
    parameter WIDTH = 8,
    parameter DEPTH = 16
)(
    input wclk,
    input rclk,
    input wrstn,
    input rrstn,
    input winc,
    input rinc,
    input [WIDTH-1:0] wdata,
    output reg wfull,
    output reg rempty,
    output reg [WIDTH-1:0] rdata
);
    localparam ADDR_WIDTH = $clog2(DEPTH);
    
    reg [ADDR_WIDTH:0] waddr_bin, raddr_bin;
    reg [ADDR_WIDTH:0] waddr_gray, raddr_gray;
    reg [ADDR_WIDTH:0] waddr_gray_d, raddr_gray_d;

    always @(posedge wclk or negedge wrstn)
        if (!wrstn)
            waddr_bin <= 0;
        else if (winc && !wfull)
            waddr_bin <= waddr_bin + 1;

    always @(posedge rclk or negedge rrstn)
        if (!rrstn)
            raddr_bin <= 0;
        else if (rinc && !rempty)
            raddr_bin <= raddr_bin + 1;

    always @(posedge wclk or negedge wrstn)
        if (!wrstn)
            waddr_gray <= 0;
        else
            waddr_gray <= waddr_bin ^ (waddr_bin >> 1);

    always @(posedge rclk or negedge rrstn)
        if (!rrstn)
            raddr_gray <= 0;
        else
            raddr_gray <= raddr_bin ^ (raddr_bin >> 1);

    always @(posedge wclk)
        waddr_gray_d <= waddr_gray;

    always @(posedge rclk)
        raddr_gray_d <= raddr_gray;

    assign wfull = (waddr_gray_d[ADDR_WIDTH:ADDR_WIDTH-1] == ~raddr_gray[ADDR_WIDTH:ADDR_WIDTH-1]) && 
                   (waddr_gray_d[ADDR_WIDTH-2:0] == raddr_gray[ADDR_WIDTH-2:0]);

    assign rempty = (waddr_gray == raddr_gray);

    wire wenc = winc && !wfull;
    wire renc = rinc && !rempty;

    dual_port_RAM #(
        .DEPTH(DEPTH),
        .WIDTH(WIDTH)
    ) RAM (
        .wclk (wclk),
        .rclk (rclk),
        .wenc (wenc),
        .waddr (waddr_bin[ADDR_WIDTH-1:0]),
        .wdata (wdata),
        .renc (renc),
        .raddr (raddr_bin[ADDR_WIDTH-1:0]),
        .rdata (rdata)
    );
endmodule
