module	asyn_fifo #(
    parameter WIDTH = 8,
    parameter DEPTH = 16
)(
    // Input ports
    input wclk,
    input rclk,
    input wrstn,
    input rrstn,
    input winc,
    input rinc,
    input [WIDTH-1:0] wdata,

    // Output ports
    output wfull,
    output rempty,
    output [WIDTH-1:0] rdata
);

    // Local parameters
    localparam ADDR_WIDTH = $clog2(DEPTH);

    // Registers and wires
    reg [ADDR_WIDTH-1:0] waddr_bin, raddr_bin, waddr_gray, raddr_gray;
    wire [ADDR_WIDTH-1:0] waddr, raddr;
    reg wenc, renc;
    reg [WIDTH-1:0] RAM[0:DEPTH-1];

    // Dual-port RAM module
    dual_port_RAM #(.DEPTH(DEPTH), .WIDTH(WIDTH)) RAM_inst (
        .wclk(wclk), .wenc(wenc), .waddr(waddr), .wdata(wdata),
        .rclk(rclk), .renc(renc), .raddr(raddr), .rdata(rdata)
    );

    // Write pointer control
    always @(posedge wclk or negedge wrstn) begin
        if (~wrstn)
            waddr_bin <= 0;
        else if (winc && !wfull)
            waddr_bin <= waddr_bin + 1;
    end

    // Read pointer control
    always @(posedge rclk or negedge rrstn) begin
        if (~rrstn)
            raddr_bin <= 0;
        else if (rinc && !rempty)
            raddr_bin <= raddr_bin + 1;
    end

    // Gray code conversion
    always @(waddr_bin) 
        waddr_gray = waddr_bin ^ (waddr_bin >> 1);
    always @(raddr_bin) 
        raddr_gray = raddr_bin ^ (raddr_bin >> 1);

    // Pointer synchronisation
    reg [ADDR_WIDTH-1:0] waddr_syn, raddr_syn;
    always @(posedge rclk or negedge rrstn) begin
        if (~rrstn)
            waddr_syn <= 0;
        else
            waddr_syn <= waddr_gray;
    end
    always @(posedge wclk or negedge wrstn) begin
        if (~wrstn)
            raddr_syn <= 0;
        else
            raddr_syn <= raddr_gray;
    end

    // Full and empty condition calculation
    assign wfull = (waddr_gray == (~raddr_syn[ADDR_WIDTH-1:ADDR_WIDTH-2], raddr_syn[ADDR_WIDTH-3:0]));
    assign rempty = (waddr_syn == raddr_gray);

    // Write and read address
    assign waddr = waddr_bin[ADDR_WIDTH-1:0];
    assign raddr = raddr_bin[ADDR_WIDTH-1:0];

    // Write and read enable
    assign wenc = winc && !wfull;
    assign renc = rinc && !rempty;

endmodule
